../../webadmin/postgresql/config.info.sv
../../webadmin/cron/config.info.sv
../../webadmin/man/config.info.sv
../../webadmin/proc/config.info.sv
desc_sv=Filhanterare
